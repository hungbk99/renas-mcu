//////////////////////////////////////////////////////////////////////////////////
// File Name: 		inst_ahb_interface.sv
// Function:		  INST-AHB Interface for renas cpu
// Project Name:	renas mcu
// Copyright (C) 	Le Quang Hung 
// Ho Chi Minh University of Technology
// Email: 			quanghungbk1999@gmail.com  
// Ver    Date        Author    Description
// v0.0   01.04.2021  hungbk99  First Creation                    
//////////////////////////////////////////////////////////////////////////////////
